library verilog;
use verilog.vl_types.all;
entity sort_tb is
end sort_tb;
