//linear search
module search(Clk,Reset);

   input Clk;
   input Reset;

	
   reg [7:0] checkx;//searches for this in queue
   reg [7:0] checky;
	
	
   reg [7:0] state;
	
   reg [7:0] closex [0:399];
   reg [7:0] closey [0:399];
   
   //output these?
   reg [8:0] search_index; //used to iterate through reg
   reg 	    found;
	
   localparam 
     CHECK_IF_IN_CLOSED	          =	8'b00_100000,
     SEARCH_CLOSED_COMPARE        = 	8'b00_100001,
     SEARCH_CLOSED_NEXT           = 	8'b00_100010,
     SEARCH_CLOSED_DONE_FOUND  	  = 	8'b00_100011,
     SEARCH_CLOSED_DONE_NOT_FOUND =  8'b00_100100;
   
	
   always @ (posedge Clk, posedge Reset)
     begin
	if(Reset)
	  begin	
	     state <= CHECK_IF_IN_CLOSED;
	     checkx <= 8'b1;
	     checky <= 8'b1;
	     
	closex[0] <= 8'b0;
closey[0] <= 8'b0;
closex[1] <= 8'b0;
closey[1] <= 8'b0;
closex[2] <= 8'b0;
closey[2] <= 8'b0;
closex[3] <= 8'b0;
closey[3] <= 8'b0;
closex[4] <= 8'b0;
closey[4] <= 8'b0;
closex[5] <= 8'b0;
closey[5] <= 8'b0;
closex[6] <= 8'b10;
closey[6] <= 8'b10;
closex[7] <= 8'b0;
closey[7] <= 8'b0;
closex[8] <= 8'b0;
closey[8] <= 8'b0;
closex[9] <= 8'b0;
closey[9] <= 8'b0;
closex[10] <= 8'b0;
closey[10] <= 8'b0;
closex[11] <= 8'b0;
closey[11] <= 8'b0;
closex[12] <= 8'b0;
closey[12] <= 8'b0;
closex[13] <= 8'b0;
closey[13] <= 8'b0;
closex[14] <= 8'b0;
closey[14] <= 8'b0;
closex[15] <= 8'b0;
closey[15] <= 8'b0;
closex[16] <= 8'b0;
closey[16] <= 8'b0;
closex[17] <= 8'b0;
closey[17] <= 8'b0;
closex[18] <= 8'b0;
closey[18] <= 8'b0;
closex[19] <= 8'b0;
closey[19] <= 8'b0;
closex[20] <= 8'b0;
closey[20] <= 8'b0;
closex[21] <= 8'b0;
closey[21] <= 8'b0;
closex[22] <= 8'b0;
closey[22] <= 8'b0;
closex[23] <= 8'b0;
closey[23] <= 8'b0;
closex[24] <= 8'b0;
closey[24] <= 8'b0;
closex[25] <= 8'b0;
closey[25] <= 8'b0;
closex[26] <= 8'b0;
closey[26] <= 8'b0;
closex[27] <= 8'b0;
closey[27] <= 8'b0;
closex[28] <= 8'b0;
closey[28] <= 8'b0;
closex[29] <= 8'b0;
closey[29] <= 8'b0;
closex[30] <= 8'b0;
closey[30] <= 8'b0;
closex[31] <= 8'b0;
closey[31] <= 8'b0;
closex[32] <= 8'b0;
closey[32] <= 8'b0;
closex[33] <= 8'b0;
closey[33] <= 8'b0;
closex[34] <= 8'b0;
closey[34] <= 8'b0;
closex[35] <= 8'b0;
closey[35] <= 8'b0;
closex[36] <= 8'b0;
closey[36] <= 8'b0;
closex[37] <= 8'b0;
closey[37] <= 8'b0;
closex[38] <= 8'b0;
closey[38] <= 8'b0;
closex[39] <= 8'b0;
closey[39] <= 8'b0;
closex[40] <= 8'b0;
closey[40] <= 8'b0;
closex[41] <= 8'b0;
closey[41] <= 8'b0;
closex[42] <= 8'b0;
closey[42] <= 8'b0;
closex[43] <= 8'b0;
closey[43] <= 8'b0;
closex[44] <= 8'b0;
closey[44] <= 8'b0;
closex[45] <= 8'b0;
closey[45] <= 8'b0;
closex[46] <= 8'b0;
closey[46] <= 8'b0;
closex[47] <= 8'b0;
closey[47] <= 8'b0;
closex[48] <= 8'b0;
closey[48] <= 8'b0;
closex[49] <= 8'b0;
closey[49] <= 8'b0;
closex[50] <= 8'b0;
closey[50] <= 8'b0;
closex[51] <= 8'b0;
closey[51] <= 8'b0;
closex[52] <= 8'b0;
closey[52] <= 8'b0;
closex[53] <= 8'b0;
closey[53] <= 8'b0;
closex[54] <= 8'b0;
closey[54] <= 8'b0;
closex[55] <= 8'b0;
closey[55] <= 8'b0;
closex[56] <= 8'b0;
closey[56] <= 8'b0;
closex[57] <= 8'b0;
closey[57] <= 8'b0;
closex[58] <= 8'b0;
closey[58] <= 8'b0;
closex[59] <= 8'b0;
closey[59] <= 8'b0;
closex[60] <= 8'b0;
closey[60] <= 8'b0;
closex[61] <= 8'b0;
closey[61] <= 8'b0;
closex[62] <= 8'b0;
closey[62] <= 8'b0;
closex[63] <= 8'b0;
closey[63] <= 8'b0;
closex[64] <= 8'b0;
closey[64] <= 8'b0;
closex[65] <= 8'b0;
closey[65] <= 8'b0;
closex[66] <= 8'b0;
closey[66] <= 8'b0;
closex[67] <= 8'b0;
closey[67] <= 8'b0;
closex[68] <= 8'b0;
closey[68] <= 8'b0;
closex[69] <= 8'b0;
closey[69] <= 8'b0;
closex[70] <= 8'b0;
closey[70] <= 8'b0;
closex[71] <= 8'b0;
closey[71] <= 8'b0;
closex[72] <= 8'b0;
closey[72] <= 8'b0;
closex[73] <= 8'b0;
closey[73] <= 8'b0;
closex[74] <= 8'b0;
closey[74] <= 8'b0;
closex[75] <= 8'b0;
closey[75] <= 8'b0;
closex[76] <= 8'b0;
closey[76] <= 8'b0;
closex[77] <= 8'b0;
closey[77] <= 8'b0;
closex[78] <= 8'b0;
closey[78] <= 8'b0;
closex[79] <= 8'b0;
closey[79] <= 8'b0;
closex[80] <= 8'b0;
closey[80] <= 8'b0;
closex[81] <= 8'b0;
closey[81] <= 8'b0;
closex[82] <= 8'b0;
closey[82] <= 8'b0;
closex[83] <= 8'b0;
closey[83] <= 8'b0;
closex[84] <= 8'b0;
closey[84] <= 8'b0;
closex[85] <= 8'b0;
closey[85] <= 8'b0;
closex[86] <= 8'b0;
closey[86] <= 8'b0;
closex[87] <= 8'b0;
closey[87] <= 8'b0;
closex[88] <= 8'b0;
closey[88] <= 8'b0;
closex[89] <= 8'b0;
closey[89] <= 8'b0;
closex[90] <= 8'b0;
closey[90] <= 8'b0;
closex[91] <= 8'b0;
closey[91] <= 8'b0;
closex[92] <= 8'b0;
closey[92] <= 8'b0;
closex[93] <= 8'b0;
closey[93] <= 8'b0;
closex[94] <= 8'b0;
closey[94] <= 8'b0;
closex[95] <= 8'b0;
closey[95] <= 8'b0;
closex[96] <= 8'b0;
closey[96] <= 8'b0;
closex[97] <= 8'b0;
closey[97] <= 8'b0;
closex[98] <= 8'b0;
closey[98] <= 8'b0;
closex[99] <= 8'b0;
closey[99] <= 8'b0;
closex[100] <= 8'b0;
closey[100] <= 8'b0;
closex[101] <= 8'b0;
closey[101] <= 8'b0;
closex[102] <= 8'b0;
closey[102] <= 8'b0;
closex[103] <= 8'b0;
closey[103] <= 8'b0;
closex[104] <= 8'b0;
closey[104] <= 8'b0;
closex[105] <= 8'b0;
closey[105] <= 8'b0;
closex[106] <= 8'b0;
closey[106] <= 8'b0;
closex[107] <= 8'b0;
closey[107] <= 8'b0;
closex[108] <= 8'b0;
closey[108] <= 8'b0;
closex[109] <= 8'b0;
closey[109] <= 8'b0;
closex[110] <= 8'b0;
closey[110] <= 8'b0;
closex[111] <= 8'b0;
closey[111] <= 8'b0;
closex[112] <= 8'b0;
closey[112] <= 8'b0;
closex[113] <= 8'b0;
closey[113] <= 8'b0;
closex[114] <= 8'b0;
closey[114] <= 8'b0;
closex[115] <= 8'b0;
closey[115] <= 8'b0;
closex[116] <= 8'b0;
closey[116] <= 8'b0;
closex[117] <= 8'b0;
closey[117] <= 8'b0;
closex[118] <= 8'b0;
closey[118] <= 8'b0;
closex[119] <= 8'b0;
closey[119] <= 8'b0;
closex[120] <= 8'b0;
closey[120] <= 8'b0;
closex[121] <= 8'b0;
closey[121] <= 8'b0;
closex[122] <= 8'b0;
closey[122] <= 8'b0;
closex[123] <= 8'b0;
closey[123] <= 8'b0;
closex[124] <= 8'b0;
closey[124] <= 8'b0;
closex[125] <= 8'b0;
closey[125] <= 8'b0;
closex[126] <= 8'b0;
closey[126] <= 8'b0;
closex[127] <= 8'b0;
closey[127] <= 8'b0;
closex[128] <= 8'b0;
closey[128] <= 8'b0;
closex[129] <= 8'b0;
closey[129] <= 8'b0;
closex[130] <= 8'b0;
closey[130] <= 8'b0;
closex[131] <= 8'b0;
closey[131] <= 8'b0;
closex[132] <= 8'b0;
closey[132] <= 8'b0;
closex[133] <= 8'b0;
closey[133] <= 8'b0;
closex[134] <= 8'b0;
closey[134] <= 8'b0;
closex[135] <= 8'b0;
closey[135] <= 8'b0;
closex[136] <= 8'b0;
closey[136] <= 8'b0;
closex[137] <= 8'b0;
closey[137] <= 8'b0;
closex[138] <= 8'b0;
closey[138] <= 8'b0;
closex[139] <= 8'b0;
closey[139] <= 8'b0;
closex[140] <= 8'b0;
closey[140] <= 8'b0;
closex[141] <= 8'b0;
closey[141] <= 8'b0;
closex[142] <= 8'b0;
closey[142] <= 8'b0;
closex[143] <= 8'b0;
closey[143] <= 8'b0;
closex[144] <= 8'b0;
closey[144] <= 8'b0;
closex[145] <= 8'b0;
closey[145] <= 8'b0;
closex[146] <= 8'b0;
closey[146] <= 8'b0;
closex[147] <= 8'b0;
closey[147] <= 8'b0;
closex[148] <= 8'b0;
closey[148] <= 8'b0;
closex[149] <= 8'b0;
closey[149] <= 8'b0;
closex[150] <= 8'b0;
closey[150] <= 8'b0;
closex[151] <= 8'b0;
closey[151] <= 8'b0;
closex[152] <= 8'b0;
closey[152] <= 8'b0;
closex[153] <= 8'b0;
closey[153] <= 8'b0;
closex[154] <= 8'b0;
closey[154] <= 8'b0;
closex[155] <= 8'b0;
closey[155] <= 8'b0;
closex[156] <= 8'b0;
closey[156] <= 8'b0;
closex[157] <= 8'b0;
closey[157] <= 8'b0;
closex[158] <= 8'b0;
closey[158] <= 8'b0;
closex[159] <= 8'b0;
closey[159] <= 8'b0;
closex[160] <= 8'b0;
closey[160] <= 8'b0;
closex[161] <= 8'b0;
closey[161] <= 8'b0;
closex[162] <= 8'b0;
closey[162] <= 8'b0;
closex[163] <= 8'b0;
closey[163] <= 8'b0;
closex[164] <= 8'b0;
closey[164] <= 8'b0;
closex[165] <= 8'b0;
closey[165] <= 8'b0;
closex[166] <= 8'b0;
closey[166] <= 8'b0;
closex[167] <= 8'b0;
closey[167] <= 8'b0;
closex[168] <= 8'b0;
closey[168] <= 8'b0;
closex[169] <= 8'b0;
closey[169] <= 8'b0;
closex[170] <= 8'b0;
closey[170] <= 8'b0;
closex[171] <= 8'b0;
closey[171] <= 8'b0;
closex[172] <= 8'b0;
closey[172] <= 8'b0;
closex[173] <= 8'b0;
closey[173] <= 8'b0;
closex[174] <= 8'b0;
closey[174] <= 8'b0;
closex[175] <= 8'b0;
closey[175] <= 8'b0;
closex[176] <= 8'b0;
closey[176] <= 8'b0;
closex[177] <= 8'b0;
closey[177] <= 8'b0;
closex[178] <= 8'b0;
closey[178] <= 8'b0;
closex[179] <= 8'b0;
closey[179] <= 8'b0;
closex[180] <= 8'b0;
closey[180] <= 8'b0;
closex[181] <= 8'b0;
closey[181] <= 8'b0;
closex[182] <= 8'b0;
closey[182] <= 8'b0;
closex[183] <= 8'b0;
closey[183] <= 8'b0;
closex[184] <= 8'b0;
closey[184] <= 8'b0;
closex[185] <= 8'b0;
closey[185] <= 8'b0;
closex[186] <= 8'b0;
closey[186] <= 8'b0;
closex[187] <= 8'b0;
closey[187] <= 8'b0;
closex[188] <= 8'b0;
closey[188] <= 8'b0;
closex[189] <= 8'b0;
closey[189] <= 8'b0;
closex[190] <= 8'b0;
closey[190] <= 8'b0;
closex[191] <= 8'b0;
closey[191] <= 8'b0;
closex[192] <= 8'b0;
closey[192] <= 8'b0;
closex[193] <= 8'b0;
closey[193] <= 8'b0;
closex[194] <= 8'b0;
closey[194] <= 8'b0;
closex[195] <= 8'b0;
closey[195] <= 8'b0;
closex[196] <= 8'b0;
closey[196] <= 8'b0;
closex[197] <= 8'b0;
closey[197] <= 8'b0;
closex[198] <= 8'b0;
closey[198] <= 8'b0;
closex[199] <= 8'b0;
closey[199] <= 8'b0;
closex[200] <= 8'b0;
closey[200] <= 8'b0;
closex[201] <= 8'b0;
closey[201] <= 8'b0;
closex[202] <= 8'b0;
closey[202] <= 8'b0;
closex[203] <= 8'b0;
closey[203] <= 8'b0;
closex[204] <= 8'b0;
closey[204] <= 8'b0;
closex[205] <= 8'b0;
closey[205] <= 8'b0;
closex[206] <= 8'b0;
closey[206] <= 8'b0;
closex[207] <= 8'b0;
closey[207] <= 8'b0;
closex[208] <= 8'b0;
closey[208] <= 8'b0;
closex[209] <= 8'b0;
closey[209] <= 8'b0;
closex[210] <= 8'b0;
closey[210] <= 8'b0;
closex[211] <= 8'b0;
closey[211] <= 8'b0;
closex[212] <= 8'b0;
closey[212] <= 8'b0;
closex[213] <= 8'b0;
closey[213] <= 8'b0;
closex[214] <= 8'b0;
closey[214] <= 8'b0;
closex[215] <= 8'b0;
closey[215] <= 8'b0;
closex[216] <= 8'b0;
closey[216] <= 8'b0;
closex[217] <= 8'b0;
closey[217] <= 8'b0;
closex[218] <= 8'b0;
closey[218] <= 8'b0;
closex[219] <= 8'b0;
closey[219] <= 8'b0;
closex[220] <= 8'b0;
closey[220] <= 8'b0;
closex[221] <= 8'b0;
closey[221] <= 8'b0;
closex[222] <= 8'b0;
closey[222] <= 8'b0;
closex[223] <= 8'b0;
closey[223] <= 8'b0;
closex[224] <= 8'b0;
closey[224] <= 8'b0;
closex[225] <= 8'b0;
closey[225] <= 8'b0;
closex[226] <= 8'b0;
closey[226] <= 8'b0;
closex[227] <= 8'b0;
closey[227] <= 8'b0;
closex[228] <= 8'b0;
closey[228] <= 8'b0;
closex[229] <= 8'b0;
closey[229] <= 8'b0;
closex[230] <= 8'b0;
closey[230] <= 8'b0;
closex[231] <= 8'b0;
closey[231] <= 8'b0;
closex[232] <= 8'b0;
closey[232] <= 8'b0;
closex[233] <= 8'b0;
closey[233] <= 8'b0;
closex[234] <= 8'b0;
closey[234] <= 8'b0;
closex[235] <= 8'b0;
closey[235] <= 8'b0;
closex[236] <= 8'b0;
closey[236] <= 8'b0;
closex[237] <= 8'b0;
closey[237] <= 8'b0;
closex[238] <= 8'b0;
closey[238] <= 8'b0;
closex[239] <= 8'b0;
closey[239] <= 8'b0;
closex[240] <= 8'b0;
closey[240] <= 8'b0;
closex[241] <= 8'b0;
closey[241] <= 8'b0;
closex[242] <= 8'b0;
closey[242] <= 8'b0;
closex[243] <= 8'b0;
closey[243] <= 8'b0;
closex[244] <= 8'b0;
closey[244] <= 8'b0;
closex[245] <= 8'b0;
closey[245] <= 8'b0;
closex[246] <= 8'b0;
closey[246] <= 8'b0;
closex[247] <= 8'b0;
closey[247] <= 8'b0;
closex[248] <= 8'b0;
closey[248] <= 8'b0;
closex[249] <= 8'b0;
closey[249] <= 8'b0;
closex[250] <= 8'b0;
closey[250] <= 8'b0;
closex[251] <= 8'b0;
closey[251] <= 8'b0;
closex[252] <= 8'b0;
closey[252] <= 8'b0;
closex[253] <= 8'b0;
closey[253] <= 8'b0;
closex[254] <= 8'b0;
closey[254] <= 8'b0;
closex[255] <= 8'b0;
closey[255] <= 8'b0;
closex[256] <= 8'b0;
closey[256] <= 8'b0;
closex[257] <= 8'b0;
closey[257] <= 8'b0;
closex[258] <= 8'b0;
closey[258] <= 8'b0;
closex[259] <= 8'b0;
closey[259] <= 8'b0;
closex[260] <= 8'b0;
closey[260] <= 8'b0;
closex[261] <= 8'b0;
closey[261] <= 8'b0;
closex[262] <= 8'b0;
closey[262] <= 8'b0;
closex[263] <= 8'b0;
closey[263] <= 8'b0;
closex[264] <= 8'b0;
closey[264] <= 8'b0;
closex[265] <= 8'b0;
closey[265] <= 8'b0;
closex[266] <= 8'b0;
closey[266] <= 8'b0;
closex[267] <= 8'b0;
closey[267] <= 8'b0;
closex[268] <= 8'b0;
closey[268] <= 8'b0;
closex[269] <= 8'b0;
closey[269] <= 8'b0;
closex[270] <= 8'b0;
closey[270] <= 8'b0;
closex[271] <= 8'b0;
closey[271] <= 8'b0;
closex[272] <= 8'b0;
closey[272] <= 8'b0;
closex[273] <= 8'b0;
closey[273] <= 8'b0;
closex[274] <= 8'b0;
closey[274] <= 8'b0;
closex[275] <= 8'b0;
closey[275] <= 8'b0;
closex[276] <= 8'b0;
closey[276] <= 8'b0;
closex[277] <= 8'b0;
closey[277] <= 8'b0;
closex[278] <= 8'b0;
closey[278] <= 8'b0;
closex[279] <= 8'b0;
closey[279] <= 8'b0;
closex[280] <= 8'b0;
closey[280] <= 8'b0;
closex[281] <= 8'b0;
closey[281] <= 8'b0;
closex[282] <= 8'b0;
closey[282] <= 8'b0;
closex[283] <= 8'b0;
closey[283] <= 8'b0;
closex[284] <= 8'b0;
closey[284] <= 8'b0;
closex[285] <= 8'b0;
closey[285] <= 8'b0;
closex[286] <= 8'b0;
closey[286] <= 8'b0;
closex[287] <= 8'b0;
closey[287] <= 8'b0;
closex[288] <= 8'b0;
closey[288] <= 8'b0;
closex[289] <= 8'b0;
closey[289] <= 8'b0;
closex[290] <= 8'b0;
closey[290] <= 8'b0;
closex[291] <= 8'b0;
closey[291] <= 8'b0;
closex[292] <= 8'b0;
closey[292] <= 8'b0;
closex[293] <= 8'b0;
closey[293] <= 8'b0;
closex[294] <= 8'b0;
closey[294] <= 8'b0;
closex[295] <= 8'b0;
closey[295] <= 8'b0;
closex[296] <= 8'b0;
closey[296] <= 8'b0;
closex[297] <= 8'b0;
closey[297] <= 8'b0;
closex[298] <= 8'b0;
closey[298] <= 8'b0;
closex[299] <= 8'b0;
closey[299] <= 8'b0;
closex[300] <= 8'b0;
closey[300] <= 8'b0;
closex[301] <= 8'b0;
closey[301] <= 8'b0;
closex[302] <= 8'b0;
closey[302] <= 8'b0;
closex[303] <= 8'b0;
closey[303] <= 8'b0;
closex[304] <= 8'b0;
closey[304] <= 8'b0;
closex[305] <= 8'b0;
closey[305] <= 8'b0;
closex[306] <= 8'b0;
closey[306] <= 8'b0;
closex[307] <= 8'b0;
closey[307] <= 8'b0;
closex[308] <= 8'b0;
closey[308] <= 8'b0;
closex[309] <= 8'b0;
closey[309] <= 8'b0;
closex[310] <= 8'b0;
closey[310] <= 8'b0;
closex[311] <= 8'b0;
closey[311] <= 8'b0;
closex[312] <= 8'b0;
closey[312] <= 8'b0;
closex[313] <= 8'b0;
closey[313] <= 8'b0;
closex[314] <= 8'b0;
closey[314] <= 8'b0;
closex[315] <= 8'b0;
closey[315] <= 8'b0;
closex[316] <= 8'b0;
closey[316] <= 8'b0;
closex[317] <= 8'b0;
closey[317] <= 8'b0;
closex[318] <= 8'b0;
closey[318] <= 8'b0;
closex[319] <= 8'b0;
closey[319] <= 8'b0;
closex[320] <= 8'b0;
closey[320] <= 8'b0;
closex[321] <= 8'b0;
closey[321] <= 8'b0;
closex[322] <= 8'b0;
closey[322] <= 8'b0;
closex[323] <= 8'b0;
closey[323] <= 8'b0;
closex[324] <= 8'b0;
closey[324] <= 8'b0;
closex[325] <= 8'b0;
closey[325] <= 8'b0;
closex[326] <= 8'b0;
closey[326] <= 8'b0;
closex[327] <= 8'b0;
closey[327] <= 8'b0;
closex[328] <= 8'b0;
closey[328] <= 8'b0;
closex[329] <= 8'b0;
closey[329] <= 8'b0;
closex[330] <= 8'b0;
closey[330] <= 8'b0;
closex[331] <= 8'b0;
closey[331] <= 8'b0;
closex[332] <= 8'b0;
closey[332] <= 8'b0;
closex[333] <= 8'b0;
closey[333] <= 8'b0;
closex[334] <= 8'b0;
closey[334] <= 8'b0;
closex[335] <= 8'b0;
closey[335] <= 8'b0;
closex[336] <= 8'b0;
closey[336] <= 8'b0;
closex[337] <= 8'b0;
closey[337] <= 8'b0;
closex[338] <= 8'b0;
closey[338] <= 8'b0;
closex[339] <= 8'b0;
closey[339] <= 8'b0;
closex[340] <= 8'b0;
closey[340] <= 8'b0;
closex[341] <= 8'b0;
closey[341] <= 8'b0;
closex[342] <= 8'b0;
closey[342] <= 8'b0;
closex[343] <= 8'b0;
closey[343] <= 8'b0;
closex[344] <= 8'b0;
closey[344] <= 8'b0;
closex[345] <= 8'b0;
closey[345] <= 8'b0;
closex[346] <= 8'b0;
closey[346] <= 8'b0;
closex[347] <= 8'b0;
closey[347] <= 8'b0;
closex[348] <= 8'b0;
closey[348] <= 8'b0;
closex[349] <= 8'b0;
closey[349] <= 8'b0;
closex[350] <= 8'b0;
closey[350] <= 8'b0;
closex[351] <= 8'b0;
closey[351] <= 8'b0;
closex[352] <= 8'b0;
closey[352] <= 8'b0;
closex[353] <= 8'b0;
closey[353] <= 8'b0;
closex[354] <= 8'b0;
closey[354] <= 8'b0;
closex[355] <= 8'b0;
closey[355] <= 8'b0;
closex[356] <= 8'b0;
closey[356] <= 8'b0;
closex[357] <= 8'b0;
closey[357] <= 8'b0;
closex[358] <= 8'b0;
closey[358] <= 8'b0;
closex[359] <= 8'b0;
closey[359] <= 8'b0;
closex[360] <= 8'b0;
closey[360] <= 8'b0;
closex[361] <= 8'b0;
closey[361] <= 8'b0;
closex[362] <= 8'b0;
closey[362] <= 8'b0;
closex[363] <= 8'b0;
closey[363] <= 8'b0;
closex[364] <= 8'b0;
closey[364] <= 8'b0;
closex[365] <= 8'b0;
closey[365] <= 8'b0;
closex[366] <= 8'b0;
closey[366] <= 8'b0;
closex[367] <= 8'b0;
closey[367] <= 8'b0;
closex[368] <= 8'b0;
closey[368] <= 8'b0;
closex[369] <= 8'b0;
closey[369] <= 8'b0;
closex[370] <= 8'b0;
closey[370] <= 8'b0;
closex[371] <= 8'b0;
closey[371] <= 8'b0;
closex[372] <= 8'b0;
closey[372] <= 8'b0;
closex[373] <= 8'b0;
closey[373] <= 8'b0;
closex[374] <= 8'b0;
closey[374] <= 8'b0;
closex[375] <= 8'b0;
closey[375] <= 8'b0;
closex[376] <= 8'b0;
closey[376] <= 8'b0;
closex[377] <= 8'b0;
closey[377] <= 8'b0;
closex[378] <= 8'b0;
closey[378] <= 8'b0;
closex[379] <= 8'b0;
closey[379] <= 8'b0;
closex[380] <= 8'b0;
closey[380] <= 8'b0;
closex[381] <= 8'b0;
closey[381] <= 8'b0;
closex[382] <= 8'b0;
closey[382] <= 8'b0;
closex[383] <= 8'b0;
closey[383] <= 8'b0;
closex[384] <= 8'b0;
closey[384] <= 8'b0;
closex[385] <= 8'b0;
closey[385] <= 8'b0;
closex[386] <= 8'b0;
closey[386] <= 8'b0;
closex[387] <= 8'b0;
closey[387] <= 8'b0;
closex[388] <= 8'b0;
closey[388] <= 8'b0;
closex[389] <= 8'b0;
closey[389] <= 8'b0;
closex[390] <= 8'b0;
closey[390] <= 8'b0;
closex[391] <= 8'b0;
closey[391] <= 8'b0;
closex[392] <= 8'b0;
closey[392] <= 8'b0;
closex[393] <= 8'b0;
closey[393] <= 8'b0;
closex[394] <= 8'b0;
closey[394] <= 8'b0;
closex[395] <= 8'b0;
closey[395] <= 8'b0;
closex[396] <= 8'b0;
closey[396] <= 8'b0;
closex[397] <= 8'b0;
closey[397] <= 8'b0;
closex[398] <= 8'b1;
closey[398] <= 8'b1;
closex[399] <= 8'b1;
closey[399] <= 8'b1;


	  end
	
	else 
	  begin
	     case(state)
////////////////////////////////////////////////////////////////////	
	       CHECK_IF_IN_CLOSED:
		 begin 
		    $display("STATE: CHECK_IF_IN_CLOSED");
		    search_index <= 9'b0;
		    found <= 1'b0;
		    state <= SEARCH_CLOSED_COMPARE;
		 end
			
	       SEARCH_CLOSED_COMPARE:
		 begin
		   $display("STATE: SEARCH_CLOSED_COMPARE");
		    if(closex[search_index] == checkx && closey[search_index] == checky)
		      begin
			 found <= 1'b1;
			 state <= SEARCH_CLOSED_DONE_FOUND; //Go to next section
		      end
		    else
		      begin
			 search_index <= search_index + 1;
			 state <= SEARCH_CLOSED_NEXT;
		      end
		 end
	       SEARCH_CLOSED_NEXT:
<<<<<<< HEAD
	       $display("STATE: SEARCH_CLOSED_NEXT");
=======
>>>>>>> 48a8114dcec4208d7e75087badb316c1c8d584b4
		 begin
		    if(search_index == closecounter)//equals 399
		      begin
			 found <=1'b0;
			 state <= SEARCH_CLOSED_DONE_NOT_FOUND; // Not found, go to next section
		      end
		    else
		      begin
			 state <=SEARCH_CLOSED_COMPARE;
		      end
		 end // case: NEXT
			SEARCH_CLOSED_DONE_FOUND:
			begin
				//state <= NEIGHBOR_CHECK_LOOP;
<<<<<<< HEAD
				$display("STATE: SEARCH_CLOSED_DONE_FOUND");
			end
	       SEARCH_CLOSED_DONE_NOT_FOUND:
	       $display("STATE: SEARCH_CLOSED_DONE_NOT_FOUND");
	       //neighborcounter <= neighborcounter + 1;
=======
				
			end
	       SEARCH_CLOSED_DONE_NOT_FOUND:
	       
>>>>>>> 48a8114dcec4208d7e75087badb316c1c8d584b4
			
		 begin
//state <= CHECK_IF_IN_OPEN;
		 end
	     

 ////////////////////////////////////////////////////////////

	     endcase // case (state)
	       
	        	     end // else: !if(Reset)
     end // always @ (posedge Clk, posedge Reset)   
endmodule // search


