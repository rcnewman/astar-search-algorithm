//linear search
module search(Clk,Reset);

   input Clk;
   input Reset;

	
   reg [7:0] checkx;//searches for this in queue
   reg [7:0] checky;
	
	
   reg [7:0] state;
	
   reg [7:0] openx [0:399];
   reg [7:0] openy [0:399];
   
   //output these?
   reg [8:0] search_index; //used to iterate through reg
   reg 	    found;
	
   localparam 
     CHECK_IF_IN_OPEN	          =	8'b00_100000,
     SEARCH_OPEN_COMPARE        = 	8'b00_100001,
     SEARCH_OPEN_NEXT           = 	8'b00_100010,
     SEARCH_OPEN_DONE_FOUND  	  = 	8'b00_100011,
     SEARCH_OPEN_DONE_NOT_FOUND =     8'b00_100100;
   
	reg [9:0] opencounter;
   
   always @ (posedge Clk, posedge Reset)
     begin
	if(Reset)
	  begin	
	     state <= CHECK_IF_IN_OPEN;
	  end
	
	else 
	  begin
	     case(state)
////////////////////////////////////////////////////////////////////	
	       CHECK_IF_IN_OPEN:
		 begin 
		    $display("STATE: CHECK_IF_IN_OPEN");
		    search_index <= 9'b0;
		    found <= 1'b0;
		    state <= SEARCH_OPEN_COMPARE;
		 end
			
	       SEARCH_OPEN_COMPARE:
		 begin
		    $display("STATE: SEARCH_OPEN_COMPARE");
		    if(openx[search_index] == checkx && openy[search_index] == checky)
		      begin
			 found <= 1'b1;
			 state <= SEARCH_OPEN_DONE_FOUND; //Go to next section
		      end
		    else
		      begin
			 search_index <= search_index + 1;
			 state <= SEARCH_OPEN_NEXT;
		      end
		 end
	       SEARCH_OPEN_NEXT:
		 begin
		    $display("STATE: SEARCH_OPEN_NEXT");
		    if(search_index == opencounter)//equals 399
		      begin
			 found <=1'b0;
			 state <= SEARCH_OPEN_DONE_NOT_FOUND; // Not found, go to next section
		      end
		    else
		      begin
			 state <=SEARCH_OPEN_COMPARE;
		      end
		 end // case: NEXT\
			SEARCH_OPEN_DONE_FOUND:
			begin
			   $display("STATE: SEARCH_OPEN_DONE_FOUND");
				//state <= CHECK_IF_NEIGHBOR_IS_BETTER;
				
			end
	       SEARCH_OPEN_DONE_NOT_FOUND:
		 begin
		    $display("STATE: SEARCH_OPEN_DONE_NOT_FOUND");
			//state <= NEIGHBOR_IS_BETTER;
			//openx[opencounter] <= tempneighborx[neighborcounter];
			//openy[opencounter] <= tempneighbory[neighborcounter];
			//opencounter <= opencounter + 1;
		 end
	     

 ////////////////////////////////////////////////////////////

	     endcase // case (state)
	       
	        	     end // else: !if(Reset)
     end // always @ (posedge Clk, posedge Reset)   
endmodule // search


