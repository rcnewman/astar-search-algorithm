module reconstruct(Clk,Reset);
  
  input Clk;
  input Reset;
  
 
  reg [7:0]   previousNodeX0 [39:0];
  reg [7:0]   previousNodeY0 [39:0];
  reg [7:0]   previousNodeX1 [39:0];
  reg [7:0]   previousNodeY1 [39:0];
  reg [7:0]   previousNodeX2 [39:0];
  reg [7:0]   previousNodeY2 [39:0];
  reg [7:0]   previousNodeX3 [39:0];
   reg [7:0]   previousNodeY3 [39:0];
   reg [7:0]   previousNodeX4 [39:0];
   reg [7:0]   previousNodeY4 [39:0];
   reg [7:0]   previousNodeX5 [39:0];
   reg [7:0]   previousNodeY5 [39:0];
   reg [7:0]   previousNodeX6 [39:0];
   reg [7:0]   previousNodeY6 [39:0];
   reg [7:0]   previousNodeX7 [39:0];
   reg [7:0]   previousNodeY7 [39:0];
   reg [7:0]   previousNodeX8 [39:0];
   reg [7:0]   previousNodeY8 [39:0];
   reg [7:0]   previousNodeX9 [39:0];
   reg [7:0]   previousNodeY9 [39:0];
   reg [7:0]   previousNodeX10 [39:0];
   reg [7:0]   previousNodeY10 [39:0];
   reg [7:0]   previousNodeX11 [39:0];
   reg [7:0]   previousNodeY11 [39:0];
   reg [7:0]   previousNodeX12 [39:0];
   reg [7:0]   previousNodeY12 [39:0];
   reg [7:0]   previousNodeX13 [39:0];
   reg [7:0]   previousNodeY13 [39:0];
   reg [7:0]   previousNodeX14 [39:0];
   reg [7:0]   previousNodeY14 [39:0];
   reg [7:0]   previousNodeX15 [39:0];
   reg [7:0]   previousNodeY15 [39:0];
   reg [7:0]   previousNodeX16 [39:0];
   reg [7:0]   previousNodeY16 [39:0];
   reg [7:0]   previousNodeX17 [39:0];
   reg [7:0]   previousNodeY17 [39:0];
   reg [7:0]   previousNodeX18 [39:0];
   reg [7:0]   previousNodeY18 [39:0];
   reg [7:0]   previousNodeX19 [39:0];
   reg [7:0]   previousNodeY19 [39:0];
   reg [7:0]   previousNodeX20 [39:0];
   reg [7:0]   previousNodeY20 [39:0];
   reg [7:0]   previousNodeX21 [39:0];
   reg [7:0]   previousNodeY21 [39:0];
   reg [7:0]   previousNodeX22 [39:0];
   reg [7:0]   previousNodeY22 [39:0];
   reg [7:0]   previousNodeX23 [39:0];
   reg [7:0]   previousNodeY23 [39:0];
   reg [7:0]   previousNodeX24 [39:0];
   reg [7:0]   previousNodeY24 [39:0];
   reg [7:0]   previousNodeX25 [39:0];
   reg [7:0]   previousNodeY25 [39:0];
   reg [7:0]   previousNodeX26 [39:0];
   reg [7:0]   previousNodeY26 [39:0];
   reg [7:0]   previousNodeX27 [39:0];
   reg [7:0]   previousNodeY27 [39:0];
   reg [7:0]   previousNodeX28 [39:0];
   reg [7:0]   previousNodeY28 [39:0];
   reg [7:0]   previousNodeX29 [39:0];
   reg [7:0]   previousNodeY29 [39:0];
   reg [7:0]   previousNodeX30 [39:0];
   reg [7:0]   previousNodeY30 [39:0];
   reg [7:0]   previousNodeX31 [39:0];
   reg [7:0]   previousNodeY31 [39:0];
   reg [7:0]   previousNodeX32 [39:0];
   reg [7:0]   previousNodeY32 [39:0];
   reg [7:0]   previousNodeX33 [39:0];
   reg [7:0]   previousNodeY33 [39:0];
   reg [7:0]   previousNodeX34 [39:0];
   reg [7:0]   previousNodeY34 [39:0];
   reg [7:0]   previousNodeX35 [39:0];
   reg [7:0]   previousNodeY35 [39:0];
   reg [7:0]   previousNodeX36 [39:0];
   reg [7:0]   previousNodeY36 [39:0];
   reg [7:0]   previousNodeX37 [39:0];
   reg [7:0]   previousNodeY37 [39:0];
   reg [7:0]   previousNodeX38 [39:0];
   reg [7:0]   previousNodeY38 [39:0];
   reg [7:0]   previousNodeX39 [39:0];
   reg [7:0]   previousNodeY39 [39:0];
   
    reg [7:0] finished_path_x [39:0];
    reg [7:0] finished_path_y [39:0];
    reg [7:0] current_recon_x;
    reg [7:0] current_recon_y;
    
localparam
	RECONSTRUCT 			= 8'000_000_00, 	
	FIND_PREVIOUS 			= 8'000_001_00,
	CHECK_RECONSTRUCT_DONE 	= 8'000_010_00,
	DONE 		= 8'000_011_00;
	
	
	always @ (posedge Clk, posedge Reset)
		begin
	if(Reset)
		begin
			state <= RECONSTRUCT;
			current_recon_x <= 8'b0000_0000;
			current_recon_y <= 8'b0000_0000;
			finished_path_x[0] <= 8'b11111111;
finished_path_y[0] <= 8'b11111111;
finished_path_x[1] <= 8'b11111111;
finished_path_y[1] <= 8'b11111111;
finished_path_x[2] <= 8'b11111111;
finished_path_y[2] <= 8'b11111111;
finished_path_x[3] <= 8'b11111111;
finished_path_y[3] <= 8'b11111111;
finished_path_x[4] <= 8'b11111111;
finished_path_y[4] <= 8'b11111111;
finished_path_x[5] <= 8'b11111111;
finished_path_y[5] <= 8'b11111111;
finished_path_x[6] <= 8'b11111111;
finished_path_y[6] <= 8'b11111111;
finished_path_x[7] <= 8'b11111111;
finished_path_y[7] <= 8'b11111111;
finished_path_x[8] <= 8'b11111111;
finished_path_y[8] <= 8'b11111111;
finished_path_x[9] <= 8'b11111111;
finished_path_y[9] <= 8'b11111111;
finished_path_x[10] <= 8'b11111111;
finished_path_y[10] <= 8'b11111111;
finished_path_x[11] <= 8'b11111111;
finished_path_y[11] <= 8'b11111111;
finished_path_x[12] <= 8'b11111111;
finished_path_y[12] <= 8'b11111111;
finished_path_x[13] <= 8'b11111111;
finished_path_y[13] <= 8'b11111111;
finished_path_x[14] <= 8'b11111111;
finished_path_y[14] <= 8'b11111111;
finished_path_x[15] <= 8'b11111111;
finished_path_y[15] <= 8'b11111111;
finished_path_x[16] <= 8'b11111111;
finished_path_y[16] <= 8'b11111111;
finished_path_x[17] <= 8'b11111111;
finished_path_y[17] <= 8'b11111111;
finished_path_x[18] <= 8'b11111111;
finished_path_y[18] <= 8'b11111111;
finished_path_x[19] <= 8'b11111111;
finished_path_y[19] <= 8'b11111111;
finished_path_x[20] <= 8'b11111111;
finished_path_y[20] <= 8'b11111111;
finished_path_x[21] <= 8'b11111111;
finished_path_y[21] <= 8'b11111111;
finished_path_x[22] <= 8'b11111111;
finished_path_y[22] <= 8'b11111111;
finished_path_x[23] <= 8'b11111111;
finished_path_y[23] <= 8'b11111111;
finished_path_x[24] <= 8'b11111111;
finished_path_y[24] <= 8'b11111111;
finished_path_x[25] <= 8'b11111111;
finished_path_y[25] <= 8'b11111111;
finished_path_x[26] <= 8'b11111111;
finished_path_y[26] <= 8'b11111111;
finished_path_x[27] <= 8'b11111111;
finished_path_y[27] <= 8'b11111111;
finished_path_x[28] <= 8'b11111111;
finished_path_y[28] <= 8'b11111111;
finished_path_x[29] <= 8'b11111111;
finished_path_y[29] <= 8'b11111111;
finished_path_x[30] <= 8'b11111111;
finished_path_y[30] <= 8'b11111111;
finished_path_x[31] <= 8'b11111111;
finished_path_y[31] <= 8'b11111111;
finished_path_x[32] <= 8'b11111111;
finished_path_y[32] <= 8'b11111111;
finished_path_x[33] <= 8'b11111111;
finished_path_y[33] <= 8'b11111111;
finished_path_x[34] <= 8'b11111111;
finished_path_y[34] <= 8'b11111111;
finished_path_x[35] <= 8'b11111111;
finished_path_y[35] <= 8'b11111111;
finished_path_x[36] <= 8'b11111111;
finished_path_y[36] <= 8'b11111111;
finished_path_x[37] <= 8'b11111111;
finished_path_y[37] <= 8'b11111111;
finished_path_x[38] <= 8'b11111111;
finished_path_y[38] <= 8'b11111111;
finished_path_x[39] <= 8'b11111111;
finished_path_y[39] <= 8'b11111111;

			recon_counter <= 0;
		end
	else begin
	case(state)
	
	
	RECONSTRUCT:
		 begin
			$display("STATE: RECONSTRUCT");
			recon_counter <= 0;
			current_recon_x <= 8'b0000_0000;
			current_recon_y <= 8'b0000_0000;
			state <= FIND_PREVIOUS;
		 end //STATE RECONSTRUCT
		 
	FIND_PREVIOUS:
	begin
		state <= CHECK_RECONSTRUCT_DONE;
		case(current_recon_x) 
			8'b0:
begin
finished_path_x[recon_counter] <= previousNodeX0[current_recon_y];
current_recon_x <= previousNodeX0[current_recon_y];
end
8'b1:
begin
finished_path_x[recon_counter] <= previousNodeX1[current_recon_y];
current_recon_x <= previousNodeX1[current_recon_y];
end
8'b10:
begin
finished_path_x[recon_counter] <= previousNodeX2[current_recon_y];
current_recon_x <= previousNodeX2[current_recon_y];
end
8'b11:
begin
finished_path_x[recon_counter] <= previousNodeX3[current_recon_y];
current_recon_x <= previousNodeX3[current_recon_y];
end
8'b100:
begin
finished_path_x[recon_counter] <= previousNodeX4[current_recon_y];
current_recon_x <= previousNodeX4[current_recon_y];
end
8'b101:
begin
finished_path_x[recon_counter] <= previousNodeX5[current_recon_y];
current_recon_x <= previousNodeX5[current_recon_y];
end
8'b110:
begin
finished_path_x[recon_counter] <= previousNodeX6[current_recon_y];
current_recon_x <= previousNodeX6[current_recon_y];
end
8'b111:
begin
finished_path_x[recon_counter] <= previousNodeX7[current_recon_y];
current_recon_x <= previousNodeX7[current_recon_y];
end
8'b1000:
begin
finished_path_x[recon_counter] <= previousNodeX8[current_recon_y];
current_recon_x <= previousNodeX8[current_recon_y];
end
8'b1001:
begin
finished_path_x[recon_counter] <= previousNodeX9[current_recon_y];
current_recon_x <= previousNodeX9[current_recon_y];
end
8'b1010:
begin
finished_path_x[recon_counter] <= previousNodeX10[current_recon_y];
current_recon_x <= previousNodeX10[current_recon_y];
end
8'b1011:
begin
finished_path_x[recon_counter] <= previousNodeX11[current_recon_y];
current_recon_x <= previousNodeX11[current_recon_y];
end
8'b1100:
begin
finished_path_x[recon_counter] <= previousNodeX12[current_recon_y];
current_recon_x <= previousNodeX12[current_recon_y];
end
8'b1101:
begin
finished_path_x[recon_counter] <= previousNodeX13[current_recon_y];
current_recon_x <= previousNodeX13[current_recon_y];
end
8'b1110:
begin
finished_path_x[recon_counter] <= previousNodeX14[current_recon_y];
current_recon_x <= previousNodeX14[current_recon_y];
end
8'b1111:
begin
finished_path_x[recon_counter] <= previousNodeX15[current_recon_y];
current_recon_x <= previousNodeX15[current_recon_y];
end
8'b10000:
begin
finished_path_x[recon_counter] <= previousNodeX16[current_recon_y];
current_recon_x <= previousNodeX16[current_recon_y];
end
8'b10001:
begin
finished_path_x[recon_counter] <= previousNodeX17[current_recon_y];
current_recon_x <= previousNodeX17[current_recon_y];
end
8'b10010:
begin
finished_path_x[recon_counter] <= previousNodeX18[current_recon_y];
current_recon_x <= previousNodeX18[current_recon_y];
end
8'b10011:
begin
finished_path_x[recon_counter] <= previousNodeX19[current_recon_y];
current_recon_x <= previousNodeX19[current_recon_y];
end
8'b10100:
begin
finished_path_x[recon_counter] <= previousNodeX20[current_recon_y];
current_recon_x <= previousNodeX20[current_recon_y];
end
8'b10101:
begin
finished_path_x[recon_counter] <= previousNodeX21[current_recon_y];
current_recon_x <= previousNodeX21[current_recon_y];
end
8'b10110:
begin
finished_path_x[recon_counter] <= previousNodeX22[current_recon_y];
current_recon_x <= previousNodeX22[current_recon_y];
end
8'b10111:
begin
finished_path_x[recon_counter] <= previousNodeX23[current_recon_y];
current_recon_x <= previousNodeX23[current_recon_y];
end
8'b11000:
begin
finished_path_x[recon_counter] <= previousNodeX24[current_recon_y];
current_recon_x <= previousNodeX24[current_recon_y];
end
8'b11001:
begin
finished_path_x[recon_counter] <= previousNodeX25[current_recon_y];
current_recon_x <= previousNodeX25[current_recon_y];
end
8'b11010:
begin
finished_path_x[recon_counter] <= previousNodeX26[current_recon_y];
current_recon_x <= previousNodeX26[current_recon_y];
end
8'b11011:
begin
finished_path_x[recon_counter] <= previousNodeX27[current_recon_y];
current_recon_x <= previousNodeX27[current_recon_y];
end
8'b11100:
begin
finished_path_x[recon_counter] <= previousNodeX28[current_recon_y];
current_recon_x <= previousNodeX28[current_recon_y];
end
8'b11101:
begin
finished_path_x[recon_counter] <= previousNodeX29[current_recon_y];
current_recon_x <= previousNodeX29[current_recon_y];
end
8'b11110:
begin
finished_path_x[recon_counter] <= previousNodeX30[current_recon_y];
current_recon_x <= previousNodeX30[current_recon_y];
end
8'b11111:
begin
finished_path_x[recon_counter] <= previousNodeX31[current_recon_y];
current_recon_x <= previousNodeX31[current_recon_y];
end
8'b100000:
begin
finished_path_x[recon_counter] <= previousNodeX32[current_recon_y];
current_recon_x <= previousNodeX32[current_recon_y];
end
8'b100001:
begin
finished_path_x[recon_counter] <= previousNodeX33[current_recon_y];
current_recon_x <= previousNodeX33[current_recon_y];
end
8'b100010:
begin
finished_path_x[recon_counter] <= previousNodeX34[current_recon_y];
current_recon_x <= previousNodeX34[current_recon_y];
end
8'b100011:
begin
finished_path_x[recon_counter] <= previousNodeX35[current_recon_y];
current_recon_x <= previousNodeX35[current_recon_y];
end
8'b100100:
begin
finished_path_x[recon_counter] <= previousNodeX36[current_recon_y];
current_recon_x <= previousNodeX36[current_recon_y];
end
8'b100101:
begin
finished_path_x[recon_counter] <= previousNodeX37[current_recon_y];
current_recon_x <= previousNodeX37[current_recon_y];
end
8'b100110:
begin
finished_path_x[recon_counter] <= previousNodeX38[current_recon_y];
current_recon_x <= previousNodeX38[current_recon_y];
end
8'b100111:
begin
finished_path_x[recon_counter] <= previousNodeX39[current_recon_y];
current_recon_x <= previousNodeX39[current_recon_y];
end
		endcase
		case(current_recon_y)
			8'b0:
begin
finished_path_y[recon_counter] <= previousNodeY0[current_recon_x];
current_recon_y <= previousNodeY0[current_recon_x];
end
8'b1:
begin
finished_path_y[recon_counter] <= previousNodeY1[current_recon_x];
current_recon_y <= previousNodeY1[current_recon_x];
end
8'b10:
begin
finished_path_y[recon_counter] <= previousNodeY2[current_recon_x];
current_recon_y <= previousNodeY2[current_recon_x];
end
8'b11:
begin
finished_path_y[recon_counter] <= previousNodeY3[current_recon_x];
current_recon_y <= previousNodeY3[current_recon_x];
end
8'b100:
begin
finished_path_y[recon_counter] <= previousNodeY4[current_recon_x];
current_recon_y <= previousNodeY4[current_recon_x];
end
8'b101:
begin
finished_path_y[recon_counter] <= previousNodeY5[current_recon_x];
current_recon_y <= previousNodeY5[current_recon_x];
end
8'b110:
begin
finished_path_y[recon_counter] <= previousNodeY6[current_recon_x];
current_recon_y <= previousNodeY6[current_recon_x];
end
8'b111:
begin
finished_path_y[recon_counter] <= previousNodeY7[current_recon_x];
current_recon_y <= previousNodeY7[current_recon_x];
end
8'b1000:
begin
finished_path_y[recon_counter] <= previousNodeY8[current_recon_x];
current_recon_y <= previousNodeY8[current_recon_x];
end
8'b1001:
begin
finished_path_y[recon_counter] <= previousNodeY9[current_recon_x];
current_recon_y <= previousNodeY9[current_recon_x];
end
8'b1010:
begin
finished_path_y[recon_counter] <= previousNodeY10[current_recon_x];
current_recon_y <= previousNodeY10[current_recon_x];
end
8'b1011:
begin
finished_path_y[recon_counter] <= previousNodeY11[current_recon_x];
current_recon_y <= previousNodeY11[current_recon_x];
end
8'b1100:
begin
finished_path_y[recon_counter] <= previousNodeY12[current_recon_x];
current_recon_y <= previousNodeY12[current_recon_x];
end
8'b1101:
begin
finished_path_y[recon_counter] <= previousNodeY13[current_recon_x];
current_recon_y <= previousNodeY13[current_recon_x];
end
8'b1110:
begin
finished_path_y[recon_counter] <= previousNodeY14[current_recon_x];
current_recon_y <= previousNodeY14[current_recon_x];
end
8'b1111:
begin
finished_path_y[recon_counter] <= previousNodeY15[current_recon_x];
current_recon_y <= previousNodeY15[current_recon_x];
end
8'b10000:
begin
finished_path_y[recon_counter] <= previousNodeY16[current_recon_x];
current_recon_y <= previousNodeY16[current_recon_x];
end
8'b10001:
begin
finished_path_y[recon_counter] <= previousNodeY17[current_recon_x];
current_recon_y <= previousNodeY17[current_recon_x];
end
8'b10010:
begin
finished_path_y[recon_counter] <= previousNodeY18[current_recon_x];
current_recon_y <= previousNodeY18[current_recon_x];
end
8'b10011:
begin
finished_path_y[recon_counter] <= previousNodeY19[current_recon_x];
current_recon_y <= previousNodeY19[current_recon_x];
end
8'b10100:
begin
finished_path_y[recon_counter] <= previousNodeY20[current_recon_x];
current_recon_y <= previousNodeY20[current_recon_x];
end
8'b10101:
begin
finished_path_y[recon_counter] <= previousNodeY21[current_recon_x];
current_recon_y <= previousNodeY21[current_recon_x];
end
8'b10110:
begin
finished_path_y[recon_counter] <= previousNodeY22[current_recon_x];
current_recon_y <= previousNodeY22[current_recon_x];
end
8'b10111:
begin
finished_path_y[recon_counter] <= previousNodeY23[current_recon_x];
current_recon_y <= previousNodeY23[current_recon_x];
end
8'b11000:
begin
finished_path_y[recon_counter] <= previousNodeY24[current_recon_x];
current_recon_y <= previousNodeY24[current_recon_x];
end
8'b11001:
begin
finished_path_y[recon_counter] <= previousNodeY25[current_recon_x];
current_recon_y <= previousNodeY25[current_recon_x];
end
8'b11010:
begin
finished_path_y[recon_counter] <= previousNodeY26[current_recon_x];
current_recon_y <= previousNodeY26[current_recon_x];
end
8'b11011:
begin
finished_path_y[recon_counter] <= previousNodeY27[current_recon_x];
current_recon_y <= previousNodeY27[current_recon_x];
end
8'b11100:
begin
finished_path_y[recon_counter] <= previousNodeY28[current_recon_x];
current_recon_y <= previousNodeY28[current_recon_x];
end
8'b11101:
begin
finished_path_y[recon_counter] <= previousNodeY29[current_recon_x];
current_recon_y <= previousNodeY29[current_recon_x];
end
8'b11110:
begin
finished_path_y[recon_counter] <= previousNodeY30[current_recon_x];
current_recon_y <= previousNodeY30[current_recon_x];
end
8'b11111:
begin
finished_path_y[recon_counter] <= previousNodeY31[current_recon_x];
current_recon_y <= previousNodeY31[current_recon_x];
end
8'b100000:
begin
finished_path_y[recon_counter] <= previousNodeY32[current_recon_x];
current_recon_y <= previousNodeY32[current_recon_x];
end
8'b100001:
begin
finished_path_y[recon_counter] <= previousNodeY33[current_recon_x];
current_recon_y <= previousNodeY33[current_recon_x];
end
8'b100010:
begin
finished_path_y[recon_counter] <= previousNodeY34[current_recon_x];
current_recon_y <= previousNodeY34[current_recon_x];
end
8'b100011:
begin
finished_path_y[recon_counter] <= previousNodeY35[current_recon_x];
current_recon_y <= previousNodeY35[current_recon_x];
end
8'b100100:
begin
finished_path_y[recon_counter] <= previousNodeY36[current_recon_x];
current_recon_y <= previousNodeY36[current_recon_x];
end
8'b100101:
begin
finished_path_y[recon_counter] <= previousNodeY37[current_recon_x];
current_recon_y <= previousNodeY37[current_recon_x];
end
8'b100110:
begin
finished_path_y[recon_counter] <= previousNodeY38[current_recon_x];
current_recon_y <= previousNodeY38[current_recon_x];
end
8'b100111:
begin
finished_path_y[recon_counter] <= previousNodeY39[current_recon_x];
current_recon_y <= previousNodeY39[current_recon_x];
end
		endcase
	end //end FIND_PREVIOUS
	
	CHECK_RECONSTRUCT_DONE;
	begin
		if(finished_path_x[recon_counter] == 0 && finished_path_y[recon_counter] == 0)
			state <= DONE;
		else
			recon_counter <= recon_counter + 1;
			state <= FIND_PREVIOUS;
	end
	DONE:
	begin
		$display("You're done mothafucka");
	end
	