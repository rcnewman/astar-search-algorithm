module test;
hey
begin
lolol
rofl
mao
end
hey  