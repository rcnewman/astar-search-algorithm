
module sort(Clk,Reset);
  
  input Clk;
  input Reset;

  reg[15:0] temp1,temp2,temp3,temp4,temp5,temp6,total1,total2;
  reg did_swap;
  
  reg [7:0] state;

  reg [399:0] openx [7:0];//open list x cord
  reg [399:0] openy [7:0];//open list y cord

  always @ (posedge Clk, posedge Reset)
  begin

    case(state)
        if(Reset)
          begin
openx[0]= 8'11111111;
openy[0]= 8'11111111;
openx[1]= 8'11111111;
openy[1]= 8'11111111;
openx[2]= 8'11111111;
openy[2]= 8'11111111;
openx[3]= 8'11111111;
openy[3]= 8'11111111;
openx[4]= 8'11111111;
openy[4]= 8'11111111;
openx[5]= 8'11111111;
openy[5]= 8'11111111;
openx[6]= 8'11111111;
openy[6]= 8'11111111;
openx[7]= 8'11111111;
openy[7]= 8'11111111;
openx[8]= 8'11111111;
openy[8]= 8'11111111;
openx[9]= 8'11111111;
openy[9]= 8'11111111;
openx[10]= 8'11111111;
openy[10]= 8'11111111;
openx[11]= 8'11111111;
openy[11]= 8'11111111;
openx[12]= 8'11111111;
openy[12]= 8'11111111;
openx[13]= 8'11111111;
openy[13]= 8'11111111;
openx[14]= 8'11111111;
openy[14]= 8'11111111;
openx[15]= 8'11111111;
openy[15]= 8'11111111;
openx[16]= 8'11111111;
openy[16]= 8'11111111;
openx[17]= 8'11111111;
openy[17]= 8'11111111;
openx[18]= 8'11111111;
openy[18]= 8'11111111;
openx[19]= 8'11111111;
openy[19]= 8'11111111;
openx[20]= 8'11111111;
openy[20]= 8'11111111;
openx[21]= 8'11111111;
openy[21]= 8'11111111;
openx[22]= 8'11111111;
openy[22]= 8'11111111;
openx[23]= 8'11111111;
openy[23]= 8'11111111;
openx[24]= 8'11111111;
openy[24]= 8'11111111;
openx[25]= 8'11111111;
openy[25]= 8'11111111;
openx[26]= 8'11111111;
openy[26]= 8'11111111;
openx[27]= 8'11111111;
openy[27]= 8'11111111;
openx[28]= 8'11111111;
openy[28]= 8'11111111;
openx[29]= 8'11111111;
openy[29]= 8'11111111;
openx[30]= 8'11111111;
openy[30]= 8'11111111;
openx[31]= 8'11111111;
openy[31]= 8'11111111;
openx[32]= 8'11111111;
openy[32]= 8'11111111;
openx[33]= 8'11111111;
openy[33]= 8'11111111;
openx[34]= 8'11111111;
openy[34]= 8'11111111;
openx[35]= 8'11111111;
openy[35]= 8'11111111;
openx[36]= 8'11111111;
openy[36]= 8'11111111;
openx[37]= 8'11111111;
openy[37]= 8'11111111;
openx[38]= 8'11111111;
openy[38]= 8'11111111;
openx[39]= 8'11111111;
openy[39]= 8'11111111;
openx[40]= 8'11111111;
openy[40]= 8'11111111;
openx[41]= 8'11111111;
openy[41]= 8'11111111;
openx[42]= 8'11111111;
openy[42]= 8'11111111;
openx[43]= 8'11111111;
openy[43]= 8'11111111;
openx[44]= 8'11111111;
openy[44]= 8'11111111;
openx[45]= 8'11111111;
openy[45]= 8'11111111;
openx[46]= 8'11111111;
openy[46]= 8'11111111;
openx[47]= 8'11111111;
openy[47]= 8'11111111;
openx[48]= 8'11111111;
openy[48]= 8'11111111;
openx[49]= 8'11111111;
openy[49]= 8'11111111;
openx[50]= 8'11111111;
openy[50]= 8'11111111;
openx[51]= 8'11111111;
openy[51]= 8'11111111;
openx[52]= 8'11111111;
openy[52]= 8'11111111;
openx[53]= 8'11111111;
openy[53]= 8'11111111;
openx[54]= 8'11111111;
openy[54]= 8'11111111;
openx[55]= 8'11111111;
openy[55]= 8'11111111;
openx[56]= 8'11111111;
openy[56]= 8'11111111;
openx[57]= 8'11111111;
openy[57]= 8'11111111;
openx[58]= 8'11111111;
openy[58]= 8'11111111;
openx[59]= 8'11111111;
openy[59]= 8'11111111;
openx[60]= 8'11111111;
openy[60]= 8'11111111;
openx[61]= 8'11111111;
openy[61]= 8'11111111;
openx[62]= 8'11111111;
openy[62]= 8'11111111;
openx[63]= 8'11111111;
openy[63]= 8'11111111;
openx[64]= 8'11111111;
openy[64]= 8'11111111;
openx[65]= 8'11111111;
openy[65]= 8'11111111;
openx[66]= 8'11111111;
openy[66]= 8'11111111;
openx[67]= 8'11111111;
openy[67]= 8'11111111;
openx[68]= 8'11111111;
openy[68]= 8'11111111;
openx[69]= 8'11111111;
openy[69]= 8'11111111;
openx[70]= 8'11111111;
openy[70]= 8'11111111;
openx[71]= 8'11111111;
openy[71]= 8'11111111;
openx[72]= 8'11111111;
openy[72]= 8'11111111;
openx[73]= 8'11111111;
openy[73]= 8'11111111;
openx[74]= 8'11111111;
openy[74]= 8'11111111;
openx[75]= 8'11111111;
openy[75]= 8'11111111;
openx[76]= 8'11111111;
openy[76]= 8'11111111;
openx[77]= 8'11111111;
openy[77]= 8'11111111;
openx[78]= 8'11111111;
openy[78]= 8'11111111;
openx[79]= 8'11111111;
openy[79]= 8'11111111;
openx[80]= 8'11111111;
openy[80]= 8'11111111;
openx[81]= 8'11111111;
openy[81]= 8'11111111;
openx[82]= 8'11111111;
openy[82]= 8'11111111;
openx[83]= 8'11111111;
openy[83]= 8'11111111;
openx[84]= 8'11111111;
openy[84]= 8'11111111;
openx[85]= 8'11111111;
openy[85]= 8'11111111;
openx[86]= 8'11111111;
openy[86]= 8'11111111;
openx[87]= 8'11111111;
openy[87]= 8'11111111;
openx[88]= 8'11111111;
openy[88]= 8'11111111;
openx[89]= 8'11111111;
openy[89]= 8'11111111;
openx[90]= 8'11111111;
openy[90]= 8'11111111;
openx[91]= 8'11111111;
openy[91]= 8'11111111;
openx[92]= 8'11111111;
openy[92]= 8'11111111;
openx[93]= 8'11111111;
openy[93]= 8'11111111;
openx[94]= 8'11111111;
openy[94]= 8'11111111;
openx[95]= 8'11111111;
openy[95]= 8'11111111;
openx[96]= 8'11111111;
openy[96]= 8'11111111;
openx[97]= 8'11111111;
openy[97]= 8'11111111;
openx[98]= 8'11111111;
openy[98]= 8'11111111;
openx[99]= 8'11111111;
openy[99]= 8'11111111;
openx[100]= 8'11111111;
openy[100]= 8'11111111;
openx[101]= 8'11111111;
openy[101]= 8'11111111;
openx[102]= 8'11111111;
openy[102]= 8'11111111;
openx[103]= 8'11111111;
openy[103]= 8'11111111;
openx[104]= 8'11111111;
openy[104]= 8'11111111;
openx[105]= 8'11111111;
openy[105]= 8'11111111;
openx[106]= 8'11111111;
openy[106]= 8'11111111;
openx[107]= 8'11111111;
openy[107]= 8'11111111;
openx[108]= 8'11111111;
openy[108]= 8'11111111;
openx[109]= 8'11111111;
openy[109]= 8'11111111;
openx[110]= 8'11111111;
openy[110]= 8'11111111;
openx[111]= 8'11111111;
openy[111]= 8'11111111;
openx[112]= 8'11111111;
openy[112]= 8'11111111;
openx[113]= 8'11111111;
openy[113]= 8'11111111;
openx[114]= 8'11111111;
openy[114]= 8'11111111;
openx[115]= 8'11111111;
openy[115]= 8'11111111;
openx[116]= 8'11111111;
openy[116]= 8'11111111;
openx[117]= 8'11111111;
openy[117]= 8'11111111;
openx[118]= 8'11111111;
openy[118]= 8'11111111;
openx[119]= 8'11111111;
openy[119]= 8'11111111;
openx[120]= 8'11111111;
openy[120]= 8'11111111;
openx[121]= 8'11111111;
openy[121]= 8'11111111;
openx[122]= 8'11111111;
openy[122]= 8'11111111;
openx[123]= 8'11111111;
openy[123]= 8'11111111;
openx[124]= 8'11111111;
openy[124]= 8'11111111;
openx[125]= 8'11111111;
openy[125]= 8'11111111;
openx[126]= 8'11111111;
openy[126]= 8'11111111;
openx[127]= 8'11111111;
openy[127]= 8'11111111;
openx[128]= 8'11111111;
openy[128]= 8'11111111;
openx[129]= 8'11111111;
openy[129]= 8'11111111;
openx[130]= 8'11111111;
openy[130]= 8'11111111;
openx[131]= 8'11111111;
openy[131]= 8'11111111;
openx[132]= 8'11111111;
openy[132]= 8'11111111;
openx[133]= 8'11111111;
openy[133]= 8'11111111;
openx[134]= 8'11111111;
openy[134]= 8'11111111;
openx[135]= 8'11111111;
openy[135]= 8'11111111;
openx[136]= 8'11111111;
openy[136]= 8'11111111;
openx[137]= 8'11111111;
openy[137]= 8'11111111;
openx[138]= 8'11111111;
openy[138]= 8'11111111;
openx[139]= 8'11111111;
openy[139]= 8'11111111;
openx[140]= 8'11111111;
openy[140]= 8'11111111;
openx[141]= 8'11111111;
openy[141]= 8'11111111;
openx[142]= 8'11111111;
openy[142]= 8'11111111;
openx[143]= 8'11111111;
openy[143]= 8'11111111;
openx[144]= 8'11111111;
openy[144]= 8'11111111;
openx[145]= 8'11111111;
openy[145]= 8'11111111;
openx[146]= 8'11111111;
openy[146]= 8'11111111;
openx[147]= 8'11111111;
openy[147]= 8'11111111;
openx[148]= 8'11111111;
openy[148]= 8'11111111;
openx[149]= 8'11111111;
openy[149]= 8'11111111;
openx[150]= 8'11111111;
openy[150]= 8'11111111;
openx[151]= 8'11111111;
openy[151]= 8'11111111;
openx[152]= 8'11111111;
openy[152]= 8'11111111;
openx[153]= 8'11111111;
openy[153]= 8'11111111;
openx[154]= 8'11111111;
openy[154]= 8'11111111;
openx[155]= 8'11111111;
openy[155]= 8'11111111;
openx[156]= 8'11111111;
openy[156]= 8'11111111;
openx[157]= 8'11111111;
openy[157]= 8'11111111;
openx[158]= 8'11111111;
openy[158]= 8'11111111;
openx[159]= 8'11111111;
openy[159]= 8'11111111;
openx[160]= 8'11111111;
openy[160]= 8'11111111;
openx[161]= 8'11111111;
openy[161]= 8'11111111;
openx[162]= 8'11111111;
openy[162]= 8'11111111;
openx[163]= 8'11111111;
openy[163]= 8'11111111;
openx[164]= 8'11111111;
openy[164]= 8'11111111;
openx[165]= 8'11111111;
openy[165]= 8'11111111;
openx[166]= 8'11111111;
openy[166]= 8'11111111;
openx[167]= 8'11111111;
openy[167]= 8'11111111;
openx[168]= 8'11111111;
openy[168]= 8'11111111;
openx[169]= 8'11111111;
openy[169]= 8'11111111;
openx[170]= 8'11111111;
openy[170]= 8'11111111;
openx[171]= 8'11111111;
openy[171]= 8'11111111;
openx[172]= 8'11111111;
openy[172]= 8'11111111;
openx[173]= 8'11111111;
openy[173]= 8'11111111;
openx[174]= 8'11111111;
openy[174]= 8'11111111;
openx[175]= 8'11111111;
openy[175]= 8'11111111;
openx[176]= 8'11111111;
openy[176]= 8'11111111;
openx[177]= 8'11111111;
openy[177]= 8'11111111;
openx[178]= 8'11111111;
openy[178]= 8'11111111;
openx[179]= 8'11111111;
openy[179]= 8'11111111;
openx[180]= 8'11111111;
openy[180]= 8'11111111;
openx[181]= 8'11111111;
openy[181]= 8'11111111;
openx[182]= 8'11111111;
openy[182]= 8'11111111;
openx[183]= 8'11111111;
openy[183]= 8'11111111;
openx[184]= 8'11111111;
openy[184]= 8'11111111;
openx[185]= 8'11111111;
openy[185]= 8'11111111;
openx[186]= 8'11111111;
openy[186]= 8'11111111;
openx[187]= 8'11111111;
openy[187]= 8'11111111;
openx[188]= 8'11111111;
openy[188]= 8'11111111;
openx[189]= 8'11111111;
openy[189]= 8'11111111;
openx[190]= 8'11111111;
openy[190]= 8'11111111;
openx[191]= 8'11111111;
openy[191]= 8'11111111;
openx[192]= 8'11111111;
openy[192]= 8'11111111;
openx[193]= 8'11111111;
openy[193]= 8'11111111;
openx[194]= 8'11111111;
openy[194]= 8'11111111;
openx[195]= 8'11111111;
openy[195]= 8'11111111;
openx[196]= 8'11111111;
openy[196]= 8'11111111;
openx[197]= 8'11111111;
openy[197]= 8'11111111;
openx[198]= 8'11111111;
openy[198]= 8'11111111;
openx[199]= 8'11111111;
openy[199]= 8'11111111;
openx[200]= 8'11111111;
openy[200]= 8'11111111;
openx[201]= 8'11111111;
openy[201]= 8'11111111;
openx[202]= 8'11111111;
openy[202]= 8'11111111;
openx[203]= 8'11111111;
openy[203]= 8'11111111;
openx[204]= 8'11111111;
openy[204]= 8'11111111;
openx[205]= 8'11111111;
openy[205]= 8'11111111;
openx[206]= 8'11111111;
openy[206]= 8'11111111;
openx[207]= 8'11111111;
openy[207]= 8'11111111;
openx[208]= 8'11111111;
openy[208]= 8'11111111;
openx[209]= 8'11111111;
openy[209]= 8'11111111;
openx[210]= 8'11111111;
openy[210]= 8'11111111;
openx[211]= 8'11111111;
openy[211]= 8'11111111;
openx[212]= 8'11111111;
openy[212]= 8'11111111;
openx[213]= 8'11111111;
openy[213]= 8'11111111;
openx[214]= 8'11111111;
openy[214]= 8'11111111;
openx[215]= 8'11111111;
openy[215]= 8'11111111;
openx[216]= 8'11111111;
openy[216]= 8'11111111;
openx[217]= 8'11111111;
openy[217]= 8'11111111;
openx[218]= 8'11111111;
openy[218]= 8'11111111;
openx[219]= 8'11111111;
openy[219]= 8'11111111;
openx[220]= 8'11111111;
openy[220]= 8'11111111;
openx[221]= 8'11111111;
openy[221]= 8'11111111;
openx[222]= 8'11111111;
openy[222]= 8'11111111;
openx[223]= 8'11111111;
openy[223]= 8'11111111;
openx[224]= 8'11111111;
openy[224]= 8'11111111;
openx[225]= 8'11111111;
openy[225]= 8'11111111;
openx[226]= 8'11111111;
openy[226]= 8'11111111;
openx[227]= 8'11111111;
openy[227]= 8'11111111;
openx[228]= 8'11111111;
openy[228]= 8'11111111;
openx[229]= 8'11111111;
openy[229]= 8'11111111;
openx[230]= 8'11111111;
openy[230]= 8'11111111;
openx[231]= 8'11111111;
openy[231]= 8'11111111;
openx[232]= 8'11111111;
openy[232]= 8'11111111;
openx[233]= 8'11111111;
openy[233]= 8'11111111;
openx[234]= 8'11111111;
openy[234]= 8'11111111;
openx[235]= 8'11111111;
openy[235]= 8'11111111;
openx[236]= 8'11111111;
openy[236]= 8'11111111;
openx[237]= 8'11111111;
openy[237]= 8'11111111;
openx[238]= 8'11111111;
openy[238]= 8'11111111;
openx[239]= 8'11111111;
openy[239]= 8'11111111;
openx[240]= 8'11111111;
openy[240]= 8'11111111;
openx[241]= 8'11111111;
openy[241]= 8'11111111;
openx[242]= 8'11111111;
openy[242]= 8'11111111;
openx[243]= 8'11111111;
openy[243]= 8'11111111;
openx[244]= 8'11111111;
openy[244]= 8'11111111;
openx[245]= 8'11111111;
openy[245]= 8'11111111;
openx[246]= 8'11111111;
openy[246]= 8'11111111;
openx[247]= 8'11111111;
openy[247]= 8'11111111;
openx[248]= 8'11111111;
openy[248]= 8'11111111;
openx[249]= 8'11111111;
openy[249]= 8'11111111;
openx[250]= 8'11111111;
openy[250]= 8'11111111;
openx[251]= 8'11111111;
openy[251]= 8'11111111;
openx[252]= 8'11111111;
openy[252]= 8'11111111;
openx[253]= 8'11111111;
openy[253]= 8'11111111;
openx[254]= 8'11111111;
openy[254]= 8'11111111;
openx[255]= 8'11111111;
openy[255]= 8'11111111;
openx[256]= 8'11111111;
openy[256]= 8'11111111;
openx[257]= 8'11111111;
openy[257]= 8'11111111;
openx[258]= 8'11111111;
openy[258]= 8'11111111;
openx[259]= 8'11111111;
openy[259]= 8'11111111;
openx[260]= 8'11111111;
openy[260]= 8'11111111;
openx[261]= 8'11111111;
openy[261]= 8'11111111;
openx[262]= 8'11111111;
openy[262]= 8'11111111;
openx[263]= 8'11111111;
openy[263]= 8'11111111;
openx[264]= 8'11111111;
openy[264]= 8'11111111;
openx[265]= 8'11111111;
openy[265]= 8'11111111;
openx[266]= 8'11111111;
openy[266]= 8'11111111;
openx[267]= 8'11111111;
openy[267]= 8'11111111;
openx[268]= 8'11111111;
openy[268]= 8'11111111;
openx[269]= 8'11111111;
openy[269]= 8'11111111;
openx[270]= 8'11111111;
openy[270]= 8'11111111;
openx[271]= 8'11111111;
openy[271]= 8'11111111;
openx[272]= 8'11111111;
openy[272]= 8'11111111;
openx[273]= 8'11111111;
openy[273]= 8'11111111;
openx[274]= 8'11111111;
openy[274]= 8'11111111;
openx[275]= 8'11111111;
openy[275]= 8'11111111;
openx[276]= 8'11111111;
openy[276]= 8'11111111;
openx[277]= 8'11111111;
openy[277]= 8'11111111;
openx[278]= 8'11111111;
openy[278]= 8'11111111;
openx[279]= 8'11111111;
openy[279]= 8'11111111;
openx[280]= 8'11111111;
openy[280]= 8'11111111;
openx[281]= 8'11111111;
openy[281]= 8'11111111;
openx[282]= 8'11111111;
openy[282]= 8'11111111;
openx[283]= 8'11111111;
openy[283]= 8'11111111;
openx[284]= 8'11111111;
openy[284]= 8'11111111;
openx[285]= 8'11111111;
openy[285]= 8'11111111;
openx[286]= 8'11111111;
openy[286]= 8'11111111;
openx[287]= 8'11111111;
openy[287]= 8'11111111;
openx[288]= 8'11111111;
openy[288]= 8'11111111;
openx[289]= 8'11111111;
openy[289]= 8'11111111;
openx[290]= 8'11111111;
openy[290]= 8'11111111;
openx[291]= 8'11111111;
openy[291]= 8'11111111;
openx[292]= 8'11111111;
openy[292]= 8'11111111;
openx[293]= 8'11111111;
openy[293]= 8'11111111;
openx[294]= 8'11111111;
openy[294]= 8'11111111;
openx[295]= 8'11111111;
openy[295]= 8'11111111;
openx[296]= 8'11111111;
openy[296]= 8'11111111;
openx[297]= 8'11111111;
openy[297]= 8'11111111;
openx[298]= 8'11111111;
openy[298]= 8'11111111;
openx[299]= 8'11111111;
openy[299]= 8'11111111;
openx[300]= 8'11111111;
openy[300]= 8'11111111;
openx[301]= 8'11111111;
openy[301]= 8'11111111;
openx[302]= 8'11111111;
openy[302]= 8'11111111;
openx[303]= 8'11111111;
openy[303]= 8'11111111;
openx[304]= 8'11111111;
openy[304]= 8'11111111;
openx[305]= 8'11111111;
openy[305]= 8'11111111;
openx[306]= 8'11111111;
openy[306]= 8'11111111;
openx[307]= 8'11111111;
openy[307]= 8'11111111;
openx[308]= 8'11111111;
openy[308]= 8'11111111;
openx[309]= 8'11111111;
openy[309]= 8'11111111;
openx[310]= 8'11111111;
openy[310]= 8'11111111;
openx[311]= 8'11111111;
openy[311]= 8'11111111;
openx[312]= 8'11111111;
openy[312]= 8'11111111;
openx[313]= 8'11111111;
openy[313]= 8'11111111;
openx[314]= 8'11111111;
openy[314]= 8'11111111;
openx[315]= 8'11111111;
openy[315]= 8'11111111;
openx[316]= 8'11111111;
openy[316]= 8'11111111;
openx[317]= 8'11111111;
openy[317]= 8'11111111;
openx[318]= 8'11111111;
openy[318]= 8'11111111;
openx[319]= 8'11111111;
openy[319]= 8'11111111;
openx[320]= 8'11111111;
openy[320]= 8'11111111;
openx[321]= 8'11111111;
openy[321]= 8'11111111;
openx[322]= 8'11111111;
openy[322]= 8'11111111;
openx[323]= 8'11111111;
openy[323]= 8'11111111;
openx[324]= 8'11111111;
openy[324]= 8'11111111;
openx[325]= 8'11111111;
openy[325]= 8'11111111;
openx[326]= 8'11111111;
openy[326]= 8'11111111;
openx[327]= 8'11111111;
openy[327]= 8'11111111;
openx[328]= 8'11111111;
openy[328]= 8'11111111;
openx[329]= 8'11111111;
openy[329]= 8'11111111;
openx[330]= 8'11111111;
openy[330]= 8'11111111;
openx[331]= 8'11111111;
openy[331]= 8'11111111;
openx[332]= 8'11111111;
openy[332]= 8'11111111;
openx[333]= 8'11111111;
openy[333]= 8'11111111;
openx[334]= 8'11111111;
openy[334]= 8'11111111;
openx[335]= 8'11111111;
openy[335]= 8'11111111;
openx[336]= 8'11111111;
openy[336]= 8'11111111;
openx[337]= 8'11111111;
openy[337]= 8'11111111;
openx[338]= 8'11111111;
openy[338]= 8'11111111;
openx[339]= 8'11111111;
openy[339]= 8'11111111;
openx[340]= 8'11111111;
openy[340]= 8'11111111;
openx[341]= 8'11111111;
openy[341]= 8'11111111;
openx[342]= 8'11111111;
openy[342]= 8'11111111;
openx[343]= 8'11111111;
openy[343]= 8'11111111;
openx[344]= 8'11111111;
openy[344]= 8'11111111;
openx[345]= 8'11111111;
openy[345]= 8'11111111;
openx[346]= 8'11111111;
openy[346]= 8'11111111;
openx[347]= 8'11111111;
openy[347]= 8'11111111;
openx[348]= 8'11111111;
openy[348]= 8'11111111;
openx[349]= 8'11111111;
openy[349]= 8'11111111;
openx[350]= 8'11111111;
openy[350]= 8'11111111;
openx[351]= 8'11111111;
openy[351]= 8'11111111;
openx[352]= 8'11111111;
openy[352]= 8'11111111;
openx[353]= 8'11111111;
openy[353]= 8'11111111;
openx[354]= 8'11111111;
openy[354]= 8'11111111;
openx[355]= 8'11111111;
openy[355]= 8'11111111;
openx[356]= 8'11111111;
openy[356]= 8'11111111;
openx[357]= 8'11111111;
openy[357]= 8'11111111;
openx[358]= 8'11111111;
openy[358]= 8'11111111;
openx[359]= 8'11111111;
openy[359]= 8'11111111;
openx[360]= 8'11111111;
openy[360]= 8'11111111;
openx[361]= 8'11111111;
openy[361]= 8'11111111;
openx[362]= 8'11111111;
openy[362]= 8'11111111;
openx[363]= 8'11111111;
openy[363]= 8'11111111;
openx[364]= 8'11111111;
openy[364]= 8'11111111;
openx[365]= 8'11111111;
openy[365]= 8'11111111;
openx[366]= 8'11111111;
openy[366]= 8'11111111;
openx[367]= 8'11111111;
openy[367]= 8'11111111;
openx[368]= 8'11111111;
openy[368]= 8'11111111;
openx[369]= 8'11111111;
openy[369]= 8'11111111;
openx[370]= 8'11111111;
openy[370]= 8'11111111;
openx[371]= 8'11111111;
openy[371]= 8'11111111;
openx[372]= 8'11111111;
openy[372]= 8'11111111;
openx[373]= 8'11111111;
openy[373]= 8'11111111;
openx[374]= 8'11111111;
openy[374]= 8'11111111;
openx[375]= 8'11111111;
openy[375]= 8'11111111;
openx[376]= 8'11111111;
openy[376]= 8'11111111;
openx[377]= 8'11111111;
openy[377]= 8'11111111;
openx[378]= 8'11111111;
openy[378]= 8'11111111;
openx[379]= 8'11111111;
openy[379]= 8'11111111;
openx[380]= 8'11111111;
openy[380]= 8'11111111;
openx[381]= 8'11111111;
openy[381]= 8'11111111;
openx[382]= 8'11111111;
openy[382]= 8'11111111;
openx[383]= 8'11111111;
openy[383]= 8'11111111;
openx[384]= 8'11111111;
openy[384]= 8'11111111;
openx[385]= 8'11111111;
openy[385]= 8'11111111;
openx[386]= 8'11111111;
openy[386]= 8'11111111;
openx[387]= 8'11111111;
openy[387]= 8'11111111;
openx[388]= 8'11111111;
openy[388]= 8'11111111;
openx[389]= 8'11111111;
openy[389]= 8'11111111;
openx[390]= 8'11111111;
openy[390]= 8'11111111;
openx[391]= 8'11111111;
openy[391]= 8'11111111;
openx[392]= 8'11111111;
openy[392]= 8'11111111;
openx[393]= 8'11111111;
openy[393]= 8'11111111;
openx[394]= 8'11111111;
openy[394]= 8'11111111;
openx[395]= 8'11111111;
openy[395]= 8'11111111;
openx[396]= 8'11111111;
openy[396]= 8'11111111;
openx[397]= 8'11111111;
openy[397]= 8'11111111;
openx[398]= 8'11111111;
openy[398]= 8'11111111;
openx[399]= 8'11111111;
openy[399]= 8'11111111;

          end
        else begin
        /////////////////////////////////////////////////////////////////////////////////
        
        
//GET FIRST, DISTANCE
BUBBLE_SORT:
	begin
	temp1 <=((openx[sort_count] - goalx < openy[sort_count] - goaly)?openy[sort_count]-goaly:openx[sort_count]-goalx);
	temp2 <= ((openy[sort_count] - goaly < 0)? -1*(openy[sort_count]-goaly):openy[sort_count]-goaly) + ((openx[sort_count]-goalx < 0)? -1 *(openx[sort_count]-goalx):openx[sort_count]-goalx);
	
	temp3 <= 1.41421 * temp1 + (temp2 - 2 * temp1);
	
	temp4 <=((openx[sort_count] - startx < openy[sort_count] - starty)?openy[sort_count]-starty:openx[sort_count]-startx);
	temp5 <= ((openy[sort_count] - starty < 0)? -1*(openy[sort_count]-starty):openy[sort_count]-starty) + ((openx[sort_count]-startx < 0)? -1 *(openx[sort_count]-startx):openx[sort_count]-startx);
	
	temp6 <= 1.41421 * temp4 + (temp5 - 2 * temp6);
	
	//TotalDistanceFromGoal
	total1 = temp3 + temp6;
	state = GET_SECOND_DISTANCE;
	end
GET_SECOND_DISTANCE:
	begin
	temp1 <=((openx[sort_count+1] - goalx < openy[sort_count+1] - goaly)?openy[sort_count+1]-goaly:openx[sort_count+1]-goalx);
	temp2 <= ((openy[sort_count+1] - goaly < 0)? -1*(openy[sort_count+1]-goaly):openy[sort_count+1]-goaly) + ((openx[sort_count+1]-goalx < 0)? -1 *(openx[sort_count+1]-goalx):openx[sort_count+1]-goalx);
	
	temp3 <= 1.41421 * temp1 + (temp2 - 2 * temp1);
	
	temp4 <=((openx[sort_count] - startx < openy[sort_count] - starty)?openy[sort_count]-starty:openx[sort_count]-startx);
	temp5 <= ((openy[sort_count+1] - starty < 0)? -1*(openy[sort_count+1]-starty):openy[sort_count+1]-starty) + ((openx[sort_count+1]-startx < 0)? -1 *(openx[sort_count+1]-startx):openx[sort_count+1]-startx);
	
	temp6 <= 1.41421 * temp4 + (temp5 - 2 * temp6);
	
	total2 = temp3 + temp6;
	end

COMPARE_BETTER:
	begin
		if(total2 > total1)
			state <= SWITCH;
		if(total1 < total2)
			state <= BUBBLE_NEXT;
	end
SWITCH:
	begin
		did_swap <= 1'b1;
		temp1 = openx[sort_count];
		openx[sort_count] = openx[sort_count+1];
		openx[sort_count+1] = sort_count;
		state <= BUBBLE_NEXT;
	end
BUBBLE_NEXT:
	begin
		if(sort_count >= open_counter && did_swap == 1'b1)
		begin
			sort_count <= 0;
			did_swap <= 1'b0;
			state <= BUBBLE_SORT;
		end
		if(sort_count >= open_counter && did_swap == 1'b0)
		begin
			sort_count <= 0;
			state <= SORT_DONE;
		end
		if(sort_count < open_counter)
		begin
			sort_count <= sort_count + 1;
			state <= BUBBLE_SORT;
		end
	end
	
	///////////////////////////////////////////////////////////////////////////
	 end
	end
endmodule;
			