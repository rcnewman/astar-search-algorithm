/*questions
 VGA output?
 string output to some sort of console for debugging? display
 */

module astar_algorithm(sync,reset,gridx,gridy,draw_grid,draw_obstacle,draw_path,draw_unknown);
   

   reg[15:0] temp1, temp2, temp3, temp4, temp5, temp6, total1, total2;//temporary calculation registers
   reg did_swap;

   reg [400] openx [7:0];//open list x cord
   reg [400] openy [7:0];//open list y cord
   reg [9]   opencounter;//count openx/y reg
   reg [400] closex [7:0];//close list x cord
   reg [400] closey [7:0];//close list y cord
   reg [9]   closecounter;//count closex/y reg

   reg [7:0] currentx;
   reg [7:0] currenty;
      
   reg 	     state[7:0];//current state
   reg 	     nextstate[7:0];//for utility sms this lets it know where to go next

   reg 	     bad;

   localparam
     INITIALIZE=8'b00000000,
     INITIALIZE_ARRAY=8'b00000001,
     VERIFY=8'b00000010,
     CHECK_DONE=8'b00000011,
     QUEUE_MODS=8'b00000100,
     SORT_QUEUE=8'b00001000,
     CREATE_NEIGHBORS=8'b00010000,
     CHECK_IF_IN_OPEN=8'b01000000,
     CHECK_IF_NEIGHBOR_IS_BETTER=8'b01100000,
     IS_BETTER=8'b01110000,
     RECONSTRUCT=8'b10000000,
     DONE=8'b11111100,
     ERROR=8'b11111111;

   reg [40]  map [39:0];
   
   always @ (posedge sync,posedge reset)
     begin
	if(reset)
	  begin
	     state <= INITIALIZE;
	  end
	else
	  begin
	case(state)
	  INITIALIZE:
	    begin
	       //STATE TRANSITION
	       state <= INITIALIZE_ARRAY;
	       //RTL
	       map[0]={0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	       map[1]={0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	       map[2]={0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	       map[3]={0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	       map[4]={0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	       map[5]={0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	       map[6]={0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	       map[7]={0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	       map[8]={0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	       map[9]={0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	       map[10]={0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	       map[11]={0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	       map[12]={0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	       map[13]={0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	       map[14]={0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	       map[15]={0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	       map[16]={0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	       map[17]={0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	       map[18]={0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	       map[19]={0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	       map[20]={0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	       map[21]={0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	       map[22]={0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	       map[23]={0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	       map[24]={0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	       map[25]={0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	       map[26]={0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	       map[27]={0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	       map[28]={0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	       map[29]={0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	       map[30]={0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	       map[31]={0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	       map[32]={0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	       map[33]={0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	       map[34]={0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	       map[35]={0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	       map[36]={0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	       map[37]={0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	       map[38]={0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	       map[39]={0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0};
	       bad = 0;
	       opencounter <= 9'b000000000;
	       closecounter <= 9'b000000000;
	       temp1 <= 32'b00000000000000000000000000000000;
	    end // case: INITIALIZE
	  INITIALIZE_ARRAY:
	    begin
	       //STATE TRANSITION
	       if(temp1 == 16'b0000000110001111)
		 state <= VERIFY;

	       //RTL
	       openx[temp1] <= 8'b11111111;
	       openy[temp1] <= 8'b11111111;
	       closex[temp1] <= 8'b11111111;
	       closey[temp1] <= 8'b11111111;
	       temp1 <= temp1 + temp1;
	    end // case: INITIALIZE_ARRAY
	  VERIFY:
	    begin
	       //TRANSITION LOGIC
	       if(map[0] == 40'b0000000000000000000000000000000000000001)
		 state <= ERROR;
	       else if(map[39] == 40'b1000000000000000000000000000000000000000)
		 state <= ERROR;
	       else
		 state <= CHECK_DONE;
	       //RTL
	       openx[0] <= 8'b00000000;
	       openy[0] <= 8'b00000000;
	       opencounter <= opencounter + 1;
	    end // case: VERIFY
	  CHECK_DONE:
	    begin
	       if(openx[0] == 8'b00100111 && openy[0] == 8'b00100111)
		 state <= RECONSTRUCT;
	       else if(openx[0] == 8'b11111111 && openy[0] == 8'b11111111)
		 state <= RECONSTRUCT;
	       else state <= QUEUE_MODS;
	    end // case: CHECK_DONE
	  QUEUE_MODS:
	    begin
	       //STATE TRANSITION
	       state <= QUEUE_MODS_SHIFT;
	       //RTL
	       currentx <= openx[0];
	       currenty <= openy[0];
	       closex[closecounter] <= openx[0];
	       closex[closecounter] <= openy[0];
	       closecounter <= closecounter + 1;
	       temp1 <= 0; 
	    end // case: QUEUE_MODS
	  QUEUE_MODS_SHIFT:
	    begin
	       //STATE TRANSITION
	       if(temp1 == 16'b0000000110001110)//equals to 398
		 state <= QUEUE_MODS_APPEND;
	       //RTL
	       openx[temp] <= openx[temp+1];
	       openy[temp] <= openy[temp+1];
	    end // case: QUEUE_MODS_SHIFT
	  QUEUE_MODS_APPEND:
	    begin
	       //STATE TRANSITION
	       state <= SORT_QUEUE;
	       //RTL
	       openx[399] <= 8'b11111111;
	       openy[399] <= 8'b11111111;
	    end // case: QUEUE_MODS_APPEND
	end // else: !if(reset)
     end // always @ (posedge sync,posedge reset)
   

   
while(openx[0] != 8'b11111111 && openy[0] != 8'b11111111)
  begin
if(openx[0] == 8'b00100111 && openy[0] == 8'b00100111)
  reconstructPath();
else
  begin
     closex[closecounter] <= openx[0];
     closey[closecounter] <= openy[0];
     closecounter <= closecounter + 1;
     popOpen();

     
     setNeighborNodes();
     for(0-numNeighbors)
       begin
if(close
       end
     
  end
     

  end





subroutine estimateDistanceToGoal(startx starty goalx goaly)
  temp1 <= ((starty-goaly < startx-goalx)?starty-goaly:startx-goalx);//h_diagonal
	    temp2 <= ((starty-goaly < 0)? -1*(starty-goaly):stary-goaly) + ((startx-goalx < 0)? -1*(startx-goalx):startx-goalx);//h_straight
	    
temp3 = 1.41421 * temp1 + (temp2 - 2*temp1);

/*
  		float h_diagonal = (float) Math.min(Math.abs(start.x-goal.x), Math.abs(start.y-goal.y));
		float h_straight = (float) (Math.abs(start.x-goal.x) + Math.abs(start.y-goal.y));
		float h_result = (float) (Math.sqrt(2) * h_diagonal + (h_straight - 2*h_diagonal));*/

   endmodule;